`define ADDITION       4'b0000
`define SUBTRACTION     4'b1000
`define AND             4'b0111
`define OR              4'b0110
`define XOR             4'b0100
`define SHIFT_LEFT      4'b0001
`define SHIFT_RIGHT     4'b0101
`define LT              4'b0010