`define LUI         7'b0110111

`define IMM_REG_ALU 7'b0010011

`define REG_REG_ALU 7'b0110011

`define LOAD        7'b0000011

`define STORE       7'b0100011

`define BRANCH      7'b1100011

`define JAL         7'b1101111

`define JALR        7'b1100111

`define AUIPC       7'b0010111