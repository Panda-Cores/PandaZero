`define LUI 7'b0110111

`define IMM_REG_ALU 7'b0010011

`define REG_REG_ALU 7'b0110011
