`define ADDITION       4'b0000
`define SHIFT_LEFT      4'b0001
`define SLT             4'b0010
`define SLTU            4'b0011
`define XOR             4'b0100
`define LSHIFT_RIGHT    4'b0101
`define OR              4'b0110
`define AND             4'b0111
`define SUBTRACTION     4'b1000
`define ASHIFT_RIGHT    4'b1101
