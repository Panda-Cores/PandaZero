`define ALU 3'b000
`define LOAD 3'b001
`define STORE 3'b001
